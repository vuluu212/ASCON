`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/26/2023 04:27:37 PM
// Design Name: 
// Module Name: s_box
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// LuT
module s_box(
    input [4:0] x,
    output reg [4:0] y
    );
    
    always @(*)
        case (x)
		5'd0: y = 5'd4;
		5'd1: y = 5'd11;
		5'd2: y = 5'd31;
		5'd3: y = 5'd20;
		5'd4: y = 5'd26;
		5'd5: y = 5'd21;
		5'd6: y = 5'd9;
		5'd7: y = 5'd2;
		5'd8: y = 5'd27;
		5'd9: y = 5'd5;
		5'd10: y = 5'd8;
		5'd11: y = 5'd18;
		5'd12: y = 5'd29;
		5'd13: y = 5'd3;
		5'd14: y = 5'd6;
		5'd15: y = 5'd28;
		5'd16: y = 5'd30;
		5'd17: y = 5'd19;
		5'd18: y = 5'd7;
		5'd19: y = 5'd14;
		5'd20: y = 5'd0;
		5'd21: y = 5'd13;
		5'd22: y = 5'd17;
		5'd23: y = 5'd24;
		5'd24: y = 5'd16;
		5'd25: y = 5'd12;
		5'd26: y = 5'd1;
		5'd27: y = 5'd25;
		5'd28: y = 5'd22;
		5'd29: y = 5'd10;
		5'd30: y = 5'd15;
		5'd31: y = 5'd23;

        default: y = 5'd0;
    endcase
endmodule


//ANF

//module s_box(input [4:0] x, output reg [4:0] y);
//    always @(x)
//    begin
//    	y[0] <= (x[0] & x[3]) ^ (x[0]) ^ (x[1]) ^ (x[3] & x[4]) ^ (x[3]);
//		y[1] <= (x[0] & x[4]) ^ (x[0]) ^ (x[1] & x[4]) ^ (x[1]) ^ (x[2]) ^ (x[3]) ^ (x[4]);
//		y[2] <= (x[0] & x[1]) ^ (x[0]) ^ (x[2]) ^ (x[3]) ^ (1);
//		y[3] <= (x[0]) ^ (x[1] & x[2]) ^ (x[1] & x[3]) ^ (x[1]) ^ (x[2] & x[3]) ^ (x[2]) ^ (x[3]) ^ (x[4]);
//		y[4] <= (x[0] & x[3]) ^ (x[1]) ^ (x[2] & x[3]) ^ (x[2]) ^ (x[3] & x[4]) ^ (x[3]) ^ (x[4]);
//	end
//endmodule



// KMAP
//module s_box(input [4:0] x, output [4:0] y);
//begin
//	assign y[0] = (x[4] & x[3] & x[1]) | (!x[4] & x[3] & !x[1]) | (!x[3] & !x[1] & x[0]) | (!x[3] & x[1] & !x[0]);
//	assign y[1] = (x[4] & x[3] & x[2]) | (x[4] & !x[3] & !x[2]) | (x[3] & x[2] & !x[1] & x[0]) | (!x[3] & !x[2] & !x[1] & x[0]) | (x[3] & x[2] & x[1] & !x[0]) | (!x[3] & !x[2] & x[1] & !x[0]) | (!x[4] & !x[3] & x[2] & x[1] & x[0]) | (!x[4] & x[3] & !x[2] & x[1] & x[0]) | (!x[4] & !x[3] & x[2] & !x[1] & !x[0]) | (!x[4] & x[3] & !x[2] & !x[1] & !x[0]);
//	assign y[2] = (x[3] & x[2] & x[1]) | (!x[3] & !x[2] & x[1]) | (x[3] & x[2] & !x[0]) | (!x[3] & !x[2] & !x[0]) | (!x[3] & x[2] & !x[1] & x[0]) | (x[3] & !x[2] & !x[1] & x[0]);
//	assign y[3] = (!x[4] & x[3] & x[2] & x[1] & x[0]) | (!x[4] & !x[3] & !x[2] & !x[1] & x[0]) | (x[4] & x[3] & x[2] & x[1] & !x[0]) | (x[4] & !x[3] & !x[2] & !x[1] & !x[0]) | (x[4] & !x[3] & x[2] & x[0]) | (x[4] & !x[2] & x[1] & x[0]) | (x[4] & x[3] & !x[1] & x[0]) | (!x[4] & !x[3] & x[2] & !x[0]) | (!x[4] & !x[2] & x[1] & !x[0]) | (!x[4] & x[3] & !x[1] & !x[0]);
//	assign y[4] = (x[3] & x[1] & x[0]) | (x[3] & !x[1] & !x[0]) | (x[4] & !x[3] & x[2] & x[1]) | (!x[4] & !x[3] & !x[2] & x[1]) | (!x[4] & !x[3] & x[2] & !x[1]) | (x[4] & !x[3] & !x[2] & !x[1]);
//end
//endmodule